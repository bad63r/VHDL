bad63r@bad63r-comp.2208:1519663835