`ifndef TEST_LIB_SV
 `define TEST_LIB_SV

`include "tests/test_base.sv"
`include "tests/test_simple.sv"

`endif
