`ifndef ALU_VERIF_PKG_SV
 `define ALU_VERIF_PKG_SV

package alu_verif_pkg;

   import umv_pkg::*;
 `include "uvm_macros.svh"

 `include "alu_config.sv"

 `include "alu_tx.sv"
 `include "alu_driver.sv"
 `include "alu_sequencer.sv"
 `include "alu_monitor.sv"
 `include "alu_agent.sv"

 `include "alu_env.sv"

 `include "sequences/alu_seq_lib.sv"
 `include "tests/test_lib.sv"
 


endpackage: alu_verif_pkg

   `include "alu_if.sv"

`endif
