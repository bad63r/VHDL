`ifndef ALU_SEQ_LIB_SV
 `define ALU_SEQ_LIB_SV

`include "sequences/alu_base_seq.sv"
`include "sequences/alu_simple_seq.sv"

`endif
